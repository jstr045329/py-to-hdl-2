library IEEE;
use IEEE.std_logic_1164.all;

entity rst_mgr is
        port(
                clk : in std_logic;
                por_0   : in  std_logic;
                rst_pb_0 : in std_logic;
                rst_log : in std_logic;
                rst_global_0 : out std_logic);
end rst_mgr;

architecture rst_mgr_arch of rst_mgr is
        signal my_bus : std_logic_vector(999 downto 0);
begin

process(clk)
begin
        if rising_edge(clk) then
sig_fast(0000) <= por or pushbutton;
sig_fast(0001) <= por or sig_fast(0000) or pushbutton;
sig_fast(0002) <= por or sig_fast(0001) or pushbutton;
sig_fast(0003) <= por or sig_fast(0002) or pushbutton;
sig_fast(0004) <= por or sig_fast(0003) or pushbutton;
sig_fast(0005) <= por or sig_fast(0004) or pushbutton;
sig_fast(0006) <= por or sig_fast(0005) or pushbutton;
sig_fast(0007) <= por or sig_fast(0006) or pushbutton;
sig_fast(0008) <= por or sig_fast(0007) or pushbutton;
sig_fast(0009) <= por or sig_fast(0008) or pushbutton;
sig_fast(0010) <= por or sig_fast(0009) or pushbutton;
sig_fast(0020) <= por or sig_fast(0019) or pushbutton;
sig_fast(0100) <= por or sig_fast(0099) or sig_fast(0081) or sig_fast(0019) or pushbutton;
sig_fast(0200) <= por or sig_fast(0199) or sig_fast(0181) or sig_fast(0119) or sig_fast(0001) or pushbutton;
sig_fast(0300) <= por or sig_fast(0299) or sig_fast(0281) or sig_fast(0219) or sig_fast(0101) or pushbutton;
sig_fast(0400) <= por or sig_fast(0399) or sig_fast(0381) or sig_fast(0319) or sig_fast(0201) or pushbutton;
sig_fast(0450) <= por or sig_fast(0449) or sig_fast(0431) or sig_fast(0369) or sig_fast(0251) or pushbutton;
sig_fast(0490) <= por or sig_fast(0489) or sig_fast(0471) or sig_fast(0409) or sig_fast(0291) or pushbutton;


sig_fast(0011) <= sig_fast(0002) or sig_fast(0002) or sig_fast(0004);
sig_fast(0012) <= sig_fast(0003) or sig_fast(0005) or sig_fast(0006);
sig_fast(0013) <= sig_fast(0009) or sig_fast(0010) or sig_fast(0008);
sig_fast(0014) <= sig_fast(0011) or sig_fast(0010) or sig_fast(0011);
sig_fast(0015) <= sig_fast(0014) or sig_fast(0013) or sig_fast(0014);
sig_fast(0016) <= sig_fast(0015) or sig_fast(0016) or sig_fast(0016);
sig_fast(0017) <= sig_fast(0017) or sig_fast(0018) or sig_fast(0005);
sig_fast(0018) <= sig_fast(0007) or sig_fast(0015) or sig_fast(0014);
sig_fast(0019) <= sig_fast(0004) or sig_fast(0017) or sig_fast(0007);
sig_fast(0021) <= sig_fast(0015) or sig_fast(0014) or sig_fast(0015);
sig_fast(0022) <= sig_fast(0019) or sig_fast(0013) or sig_fast(0017);
sig_fast(0023) <= sig_fast(0018) or sig_fast(0019) or sig_fast(0019);
sig_fast(0024) <= sig_fast(0020) or sig_fast(0022) or sig_fast(0018);
sig_fast(0025) <= sig_fast(0020) or sig_fast(0006) or sig_fast(0009);
sig_fast(0026) <= sig_fast(0016) or sig_fast(0003) or sig_fast(0013);
sig_fast(0027) <= sig_fast(0021) or sig_fast(0007) or sig_fast(0010);
sig_fast(0028) <= sig_fast(0009) or sig_fast(0009) or sig_fast(0015);
sig_fast(0029) <= sig_fast(0028) or sig_fast(0012) or sig_fast(0013);
sig_fast(0030) <= sig_fast(0016) or sig_fast(0023) or sig_fast(0019);
sig_fast(0031) <= sig_fast(0026) or sig_fast(0029) or sig_fast(0028);
sig_fast(0032) <= sig_fast(0001) or sig_fast(0009) or sig_fast(0027);
sig_fast(0033) <= sig_fast(0017) or sig_fast(0018) or sig_fast(0005);
sig_fast(0034) <= sig_fast(0020) or sig_fast(0014) or sig_fast(0023);
sig_fast(0035) <= sig_fast(0031) or sig_fast(0014) or sig_fast(0033);
sig_fast(0036) <= sig_fast(0019) or sig_fast(0033) or sig_fast(0019);
sig_fast(0037) <= sig_fast(0019) or sig_fast(0023) or sig_fast(0028);
sig_fast(0038) <= sig_fast(0025) or sig_fast(0020) or sig_fast(0035);
sig_fast(0039) <= sig_fast(0032) or sig_fast(0022) or sig_fast(0012);
sig_fast(0040) <= sig_fast(0036) or sig_fast(0026) or sig_fast(0006) or pushbutton;
sig_fast(0041) <= sig_fast(0032) or sig_fast(0013) or sig_fast(0031);
sig_fast(0042) <= sig_fast(0037) or sig_fast(0027) or sig_fast(0031);
sig_fast(0043) <= sig_fast(0034) or sig_fast(0019) or sig_fast(0015);
sig_fast(0044) <= sig_fast(0032) or sig_fast(0038) or sig_fast(0026);
sig_fast(0045) <= sig_fast(0026) or sig_fast(0006) or sig_fast(0006);
sig_fast(0046) <= sig_fast(0004) or sig_fast(0044) or sig_fast(0030);
sig_fast(0047) <= sig_fast(0006) or sig_fast(0019) or sig_fast(0025);
sig_fast(0048) <= sig_fast(0035) or sig_fast(0037) or sig_fast(0022);
sig_fast(0049) <= sig_fast(0020) or sig_fast(0031) or sig_fast(0014);
sig_fast(0050) <= sig_fast(0044) or sig_fast(0043) or sig_fast(0023);
sig_fast(0051) <= sig_fast(0018) or sig_fast(0018) or sig_fast(0027);
sig_fast(0052) <= sig_fast(0000) or sig_fast(0048) or sig_fast(0044);
sig_fast(0053) <= sig_fast(0045) or sig_fast(0030) or sig_fast(0033);
sig_fast(0054) <= sig_fast(0032) or sig_fast(0042) or sig_fast(0031);
sig_fast(0055) <= sig_fast(0024) or sig_fast(0016) or sig_fast(0052);
sig_fast(0056) <= sig_fast(0046) or sig_fast(0016) or sig_fast(0040);
sig_fast(0057) <= sig_fast(0038) or sig_fast(0017) or sig_fast(0050);
sig_fast(0058) <= sig_fast(0038) or sig_fast(0025) or sig_fast(0039);
sig_fast(0059) <= sig_fast(0054) or sig_fast(0025) or sig_fast(0043);
sig_fast(0060) <= sig_fast(0023) or sig_fast(0007) or sig_fast(0018) or pushbutton;
sig_fast(0061) <= sig_fast(0025) or sig_fast(0036) or sig_fast(0027);
sig_fast(0062) <= sig_fast(0017) or sig_fast(0048) or sig_fast(0039);
sig_fast(0063) <= sig_fast(0026) or sig_fast(0061) or sig_fast(0054);
sig_fast(0064) <= sig_fast(0049) or sig_fast(0060) or sig_fast(0056);
sig_fast(0065) <= sig_fast(0044) or sig_fast(0006) or sig_fast(0034);
sig_fast(0066) <= sig_fast(0021) or sig_fast(0051) or sig_fast(0040);
sig_fast(0067) <= sig_fast(0005) or sig_fast(0061) or sig_fast(0016);
sig_fast(0068) <= sig_fast(0011) or sig_fast(0057) or sig_fast(0061);
sig_fast(0069) <= sig_fast(0030) or sig_fast(0053) or sig_fast(0029);
sig_fast(0070) <= sig_fast(0069) or sig_fast(0019) or sig_fast(0028);
sig_fast(0071) <= sig_fast(0063) or sig_fast(0019) or sig_fast(0047);
sig_fast(0072) <= sig_fast(0044) or sig_fast(0024) or sig_fast(0052);
sig_fast(0073) <= sig_fast(0014) or sig_fast(0044) or sig_fast(0008);
sig_fast(0074) <= sig_fast(0044) or sig_fast(0007) or sig_fast(0042);
sig_fast(0075) <= sig_fast(0052) or sig_fast(0074) or sig_fast(0030);
sig_fast(0076) <= sig_fast(0041) or sig_fast(0064) or sig_fast(0028);
sig_fast(0077) <= sig_fast(0059) or sig_fast(0024) or sig_fast(0049);
sig_fast(0078) <= sig_fast(0069) or sig_fast(0039) or sig_fast(0026);
sig_fast(0079) <= sig_fast(0017) or sig_fast(0029) or sig_fast(0056);
sig_fast(0080) <= sig_fast(0060) or sig_fast(0038) or sig_fast(0064) or pushbutton;
sig_fast(0081) <= sig_fast(0052) or sig_fast(0046) or sig_fast(0048);
sig_fast(0082) <= sig_fast(0020) or sig_fast(0051) or sig_fast(0025);
sig_fast(0083) <= sig_fast(0060) or sig_fast(0074) or sig_fast(0017);
sig_fast(0084) <= sig_fast(0080) or sig_fast(0048) or sig_fast(0060);
sig_fast(0085) <= sig_fast(0030) or sig_fast(0026) or sig_fast(0035);
sig_fast(0086) <= sig_fast(0052) or sig_fast(0029) or sig_fast(0055);
sig_fast(0087) <= sig_fast(0054) or sig_fast(0013) or sig_fast(0080);
sig_fast(0088) <= sig_fast(0073) or sig_fast(0034) or sig_fast(0053);
sig_fast(0089) <= sig_fast(0027) or sig_fast(0053) or sig_fast(0018);
sig_fast(0090) <= sig_fast(0047) or sig_fast(0053) or sig_fast(0033);
sig_fast(0091) <= sig_fast(0022) or sig_fast(0045) or sig_fast(0086);
sig_fast(0092) <= sig_fast(0006) or sig_fast(0017) or sig_fast(0075);
sig_fast(0093) <= sig_fast(0052) or sig_fast(0045) or sig_fast(0063);
sig_fast(0094) <= sig_fast(0007) or sig_fast(0048) or sig_fast(0065);
sig_fast(0095) <= sig_fast(0045) or sig_fast(0044) or sig_fast(0093);
sig_fast(0096) <= sig_fast(0084) or sig_fast(0041) or sig_fast(0035);
sig_fast(0097) <= sig_fast(0076) or sig_fast(0039) or sig_fast(0052);
sig_fast(0098) <= sig_fast(0076) or sig_fast(0031) or sig_fast(0069);
sig_fast(0099) <= sig_fast(0028) or sig_fast(0043) or sig_fast(0062);
sig_fast(0101) <= sig_fast(0005) or sig_fast(0084) or sig_fast(0062);
sig_fast(0102) <= sig_fast(0065) or sig_fast(0019) or sig_fast(0015);
sig_fast(0103) <= sig_fast(0072) or sig_fast(0036) or sig_fast(0066);
sig_fast(0104) <= sig_fast(0066) or sig_fast(0086) or sig_fast(0020);
sig_fast(0105) <= sig_fast(0083) or sig_fast(0063) or sig_fast(0101);
sig_fast(0106) <= sig_fast(0097) or sig_fast(0014) or sig_fast(0069);
sig_fast(0107) <= sig_fast(0035) or sig_fast(0017) or sig_fast(0103);
sig_fast(0108) <= sig_fast(0028) or sig_fast(0028) or sig_fast(0094);
sig_fast(0109) <= sig_fast(0027) or sig_fast(0094) or sig_fast(0082);
sig_fast(0110) <= sig_fast(0027) or sig_fast(0040) or sig_fast(0026);
sig_fast(0111) <= sig_fast(0021) or sig_fast(0081) or sig_fast(0098);
sig_fast(0112) <= sig_fast(0076) or sig_fast(0032) or sig_fast(0044);
sig_fast(0113) <= sig_fast(0083) or sig_fast(0020) or sig_fast(0022);
sig_fast(0114) <= sig_fast(0106) or sig_fast(0076) or sig_fast(0017);
sig_fast(0115) <= sig_fast(0007) or sig_fast(0070) or sig_fast(0011);
sig_fast(0116) <= sig_fast(0018) or sig_fast(0092) or sig_fast(0082);
sig_fast(0117) <= sig_fast(0056) or sig_fast(0016) or sig_fast(0081);
sig_fast(0118) <= sig_fast(0039) or sig_fast(0021) or sig_fast(0091);
sig_fast(0119) <= sig_fast(0027) or sig_fast(0093) or sig_fast(0002);
sig_fast(0120) <= sig_fast(0013) or sig_fast(0082) or sig_fast(0014) or pushbutton;
sig_fast(0121) <= sig_fast(0033) or sig_fast(0007) or sig_fast(0076);
sig_fast(0122) <= sig_fast(0064) or sig_fast(0115) or sig_fast(0024);
sig_fast(0123) <= sig_fast(0013) or sig_fast(0120) or sig_fast(0101);
sig_fast(0124) <= sig_fast(0108) or sig_fast(0094) or sig_fast(0041);
sig_fast(0125) <= sig_fast(0105) or sig_fast(0034) or sig_fast(0044);
sig_fast(0126) <= sig_fast(0048) or sig_fast(0112) or sig_fast(0067);
sig_fast(0127) <= sig_fast(0055) or sig_fast(0091) or sig_fast(0028);
sig_fast(0128) <= sig_fast(0074) or sig_fast(0033) or sig_fast(0085);
sig_fast(0129) <= sig_fast(0066) or sig_fast(0126) or sig_fast(0014);
sig_fast(0130) <= sig_fast(0114) or sig_fast(0062) or sig_fast(0115);
sig_fast(0131) <= sig_fast(0093) or sig_fast(0129) or sig_fast(0056);
sig_fast(0132) <= sig_fast(0034) or sig_fast(0102) or sig_fast(0116);
sig_fast(0133) <= sig_fast(0056) or sig_fast(0011) or sig_fast(0047);
sig_fast(0134) <= sig_fast(0122) or sig_fast(0051) or sig_fast(0133);
sig_fast(0135) <= sig_fast(0106) or sig_fast(0044) or sig_fast(0104);
sig_fast(0136) <= sig_fast(0080) or sig_fast(0067) or sig_fast(0085);
sig_fast(0137) <= sig_fast(0060) or sig_fast(0039) or sig_fast(0061);
sig_fast(0138) <= sig_fast(0031) or sig_fast(0033) or sig_fast(0094);
sig_fast(0139) <= sig_fast(0100) or sig_fast(0137) or sig_fast(0024);
sig_fast(0140) <= sig_fast(0022) or sig_fast(0102) or sig_fast(0091) or pushbutton;
sig_fast(0141) <= sig_fast(0051) or sig_fast(0019) or sig_fast(0032);
sig_fast(0142) <= sig_fast(0046) or sig_fast(0017) or sig_fast(0121);
sig_fast(0143) <= sig_fast(0127) or sig_fast(0061) or sig_fast(0085);
sig_fast(0144) <= sig_fast(0104) or sig_fast(0135) or sig_fast(0096);
sig_fast(0145) <= sig_fast(0063) or sig_fast(0138) or sig_fast(0118);
sig_fast(0146) <= sig_fast(0045) or sig_fast(0095) or sig_fast(0143);
sig_fast(0147) <= sig_fast(0107) or sig_fast(0105) or sig_fast(0009);
sig_fast(0148) <= sig_fast(0143) or sig_fast(0130) or sig_fast(0061);
sig_fast(0149) <= sig_fast(0038) or sig_fast(0033) or sig_fast(0111);
sig_fast(0150) <= sig_fast(0084) or sig_fast(0049) or sig_fast(0036);
sig_fast(0151) <= sig_fast(0142) or sig_fast(0145) or sig_fast(0069);
sig_fast(0152) <= sig_fast(0090) or sig_fast(0032) or sig_fast(0047);
sig_fast(0153) <= sig_fast(0130) or sig_fast(0087) or sig_fast(0090);
sig_fast(0154) <= sig_fast(0026) or sig_fast(0097) or sig_fast(0153);
sig_fast(0155) <= sig_fast(0067) or sig_fast(0037) or sig_fast(0116);
sig_fast(0156) <= sig_fast(0138) or sig_fast(0032) or sig_fast(0053);
sig_fast(0157) <= sig_fast(0079) or sig_fast(0072) or sig_fast(0151);
sig_fast(0158) <= sig_fast(0091) or sig_fast(0043) or sig_fast(0051);
sig_fast(0159) <= sig_fast(0140) or sig_fast(0056) or sig_fast(0020);
sig_fast(0160) <= sig_fast(0065) or sig_fast(0002) or sig_fast(0034) or pushbutton;
sig_fast(0161) <= sig_fast(0084) or sig_fast(0135) or sig_fast(0031);
sig_fast(0162) <= sig_fast(0097) or sig_fast(0118) or sig_fast(0046);
sig_fast(0163) <= sig_fast(0156) or sig_fast(0137) or sig_fast(0115);
sig_fast(0164) <= sig_fast(0121) or sig_fast(0133) or sig_fast(0034);
sig_fast(0165) <= sig_fast(0143) or sig_fast(0040) or sig_fast(0049);
sig_fast(0166) <= sig_fast(0164) or sig_fast(0005) or sig_fast(0161);
sig_fast(0167) <= sig_fast(0059) or sig_fast(0018) or sig_fast(0042);
sig_fast(0168) <= sig_fast(0066) or sig_fast(0042) or sig_fast(0110);
sig_fast(0169) <= sig_fast(0103) or sig_fast(0101) or sig_fast(0016);
sig_fast(0170) <= sig_fast(0087) or sig_fast(0013) or sig_fast(0128);
sig_fast(0171) <= sig_fast(0151) or sig_fast(0033) or sig_fast(0094);
sig_fast(0172) <= sig_fast(0030) or sig_fast(0116) or sig_fast(0079);
sig_fast(0173) <= sig_fast(0149) or sig_fast(0085) or sig_fast(0014);
sig_fast(0174) <= sig_fast(0108) or sig_fast(0170) or sig_fast(0059);
sig_fast(0175) <= sig_fast(0100) or sig_fast(0151) or sig_fast(0169);
sig_fast(0176) <= sig_fast(0156) or sig_fast(0111) or sig_fast(0081);
sig_fast(0177) <= sig_fast(0096) or sig_fast(0055) or sig_fast(0116);
sig_fast(0178) <= sig_fast(0168) or sig_fast(0049) or sig_fast(0124);
sig_fast(0179) <= sig_fast(0024) or sig_fast(0116) or sig_fast(0140);
sig_fast(0180) <= sig_fast(0011) or sig_fast(0152) or sig_fast(0013) or pushbutton;
sig_fast(0181) <= sig_fast(0007) or sig_fast(0180) or sig_fast(0026);
sig_fast(0182) <= sig_fast(0098) or sig_fast(0042) or sig_fast(0061);
sig_fast(0183) <= sig_fast(0162) or sig_fast(0034) or sig_fast(0110);
sig_fast(0184) <= sig_fast(0141) or sig_fast(0159) or sig_fast(0151);
sig_fast(0185) <= sig_fast(0096) or sig_fast(0183) or sig_fast(0104);
sig_fast(0186) <= sig_fast(0079) or sig_fast(0009) or sig_fast(0163);
sig_fast(0187) <= sig_fast(0112) or sig_fast(0030) or sig_fast(0014);
sig_fast(0188) <= sig_fast(0046) or sig_fast(0162) or sig_fast(0096);
sig_fast(0189) <= sig_fast(0075) or sig_fast(0057) or sig_fast(0099);
sig_fast(0190) <= sig_fast(0096) or sig_fast(0167) or sig_fast(0069);
sig_fast(0191) <= sig_fast(0038) or sig_fast(0016) or sig_fast(0075);
sig_fast(0192) <= sig_fast(0103) or sig_fast(0107) or sig_fast(0161);
sig_fast(0193) <= sig_fast(0029) or sig_fast(0188) or sig_fast(0142);
sig_fast(0194) <= sig_fast(0150) or sig_fast(0039) or sig_fast(0087);
sig_fast(0195) <= sig_fast(0159) or sig_fast(0099) or sig_fast(0073);
sig_fast(0196) <= sig_fast(0096) or sig_fast(0154) or sig_fast(0077);
sig_fast(0197) <= sig_fast(0110) or sig_fast(0022) or sig_fast(0187);
sig_fast(0198) <= sig_fast(0193) or sig_fast(0071) or sig_fast(0067);
sig_fast(0199) <= sig_fast(0071) or sig_fast(0123) or sig_fast(0100);
sig_slow(0) <= sig_fast(0);
sig_slow(0001) <= sig_slow(0000) or sig_fast(0142) or sig_slow(0000) or sig_slow(0000) or sig_slow(0000);
sig_slow(0002) <= sig_slow(0001) or sig_fast(0003) or sig_slow(0000) or sig_slow(0001) or sig_slow(0000);
sig_slow(0003) <= sig_slow(0002) or sig_fast(0049) or sig_slow(0002) or sig_slow(0001) or sig_slow(0000);
sig_slow(0004) <= sig_slow(0003) or sig_fast(0074) or sig_slow(0003) or sig_slow(0003) or sig_slow(0003);
sig_slow(0005) <= sig_slow(0004) or sig_fast(0008) or sig_slow(0003) or sig_slow(0003) or sig_slow(0002);
sig_slow(0006) <= sig_slow(0005) or sig_fast(0062) or sig_slow(0001) or sig_slow(0005) or sig_slow(0005);
sig_slow(0007) <= sig_slow(0006) or sig_fast(0066) or sig_slow(0002) or sig_slow(0003) or sig_slow(0000);
sig_slow(0008) <= sig_slow(0007) or sig_fast(0132) or sig_slow(0002) or sig_slow(0007) or sig_slow(0003);
sig_slow(0009) <= sig_slow(0008) or sig_fast(0057) or sig_slow(0006) or sig_slow(0002) or sig_slow(0003);
sig_slow(0010) <= sig_slow(0009) or sig_fast(0094) or sig_slow(0007) or sig_slow(0000) or sig_slow(0003);
sig_slow(0011) <= sig_slow(0010) or sig_fast(0029) or sig_slow(0009) or sig_slow(0001) or sig_slow(0000);
sig_slow(0012) <= sig_slow(0011) or sig_fast(0085) or sig_slow(0006) or sig_slow(0001) or sig_slow(0011);
sig_slow(0013) <= sig_slow(0012) or sig_fast(0106) or sig_slow(0004) or sig_slow(0005) or sig_slow(0004);
sig_slow(0014) <= sig_slow(0013) or sig_fast(0155) or sig_slow(0008) or sig_slow(0005) or sig_slow(0007);
sig_slow(0015) <= sig_slow(0014) or sig_fast(0006) or sig_slow(0001) or sig_slow(0008) or sig_slow(0007);
sig_slow(0016) <= sig_slow(0015) or sig_fast(0062) or sig_slow(0000) or sig_slow(0002) or sig_slow(0002);
sig_slow(0017) <= sig_slow(0016) or sig_fast(0148) or sig_slow(0002) or sig_slow(0011) or sig_slow(0016);
sig_slow(0018) <= sig_slow(0017) or sig_fast(0027) or sig_slow(0014) or sig_slow(0015) or sig_slow(0003);
sig_slow(0019) <= sig_slow(0018) or sig_fast(0184) or sig_slow(0010) or sig_slow(0007) or sig_slow(0004);
sig_slow(0020) <= sig_slow(0019) or sig_fast(0128) or sig_slow(0004) or sig_slow(0005) or sig_slow(0018) or pushbutton;
sig_slow(0021) <= sig_slow(0020) or sig_fast(0146) or sig_slow(0002) or sig_slow(0014) or sig_slow(0001);
sig_slow(0022) <= sig_slow(0021) or sig_fast(0155) or sig_slow(0018) or sig_slow(0001) or sig_slow(0015);
sig_slow(0023) <= sig_slow(0022) or sig_fast(0054) or sig_slow(0015) or sig_slow(0000) or sig_slow(0012);
sig_slow(0024) <= sig_slow(0023) or sig_fast(0030) or sig_slow(0018) or sig_slow(0016) or sig_slow(0013);
sig_slow(0025) <= sig_slow(0024) or sig_fast(0184) or sig_slow(0017) or sig_slow(0012) or sig_slow(0006);
sig_slow(0026) <= sig_slow(0025) or sig_fast(0032) or sig_slow(0005) or sig_slow(0002) or sig_slow(0013);
sig_slow(0027) <= sig_slow(0026) or sig_fast(0101) or sig_slow(0025) or sig_slow(0000) or sig_slow(0009);
sig_slow(0028) <= sig_slow(0027) or sig_fast(0127) or sig_slow(0005) or sig_slow(0024) or sig_slow(0018);
sig_slow(0029) <= sig_slow(0028) or sig_fast(0094) or sig_slow(0023) or sig_slow(0008) or sig_slow(0019);
sig_slow(0030) <= sig_slow(0029) or sig_fast(0137) or sig_slow(0028) or sig_slow(0010) or sig_slow(0016);
sig_slow(0031) <= sig_slow(0030) or sig_fast(0053) or sig_slow(0014) or sig_slow(0025) or sig_slow(0000);
sig_slow(0032) <= sig_slow(0031) or sig_fast(0194) or sig_slow(0026) or sig_slow(0029) or sig_slow(0029);
sig_slow(0033) <= sig_slow(0032) or sig_fast(0037) or sig_slow(0032) or sig_slow(0012) or sig_slow(0022);
sig_slow(0034) <= sig_slow(0033) or sig_fast(0088) or sig_slow(0016) or sig_slow(0021) or sig_slow(0005);
sig_slow(0035) <= sig_slow(0034) or sig_fast(0147) or sig_slow(0017) or sig_slow(0001) or sig_slow(0016);
sig_slow(0036) <= sig_slow(0035) or sig_fast(0048) or sig_slow(0025) or sig_slow(0027) or sig_slow(0014);
sig_slow(0037) <= sig_slow(0036) or sig_fast(0026) or sig_slow(0032) or sig_slow(0009) or sig_slow(0023);
sig_slow(0038) <= sig_slow(0037) or sig_fast(0067) or sig_slow(0001) or sig_slow(0031) or sig_slow(0019);
sig_slow(0039) <= sig_slow(0038) or sig_fast(0109) or sig_slow(0022) or sig_slow(0021) or sig_slow(0009);
sig_slow(0040) <= sig_slow(0039) or sig_fast(0157) or sig_slow(0015) or sig_slow(0017) or sig_slow(0005) or pushbutton;
sig_slow(0041) <= sig_slow(0040) or sig_fast(0161) or sig_slow(0018) or sig_slow(0007) or sig_slow(0020);
sig_slow(0042) <= sig_slow(0041) or sig_fast(0034) or sig_slow(0025) or sig_slow(0016) or sig_slow(0024);
sig_slow(0043) <= sig_slow(0042) or sig_fast(0065) or sig_slow(0033) or sig_slow(0003) or sig_slow(0024);
sig_slow(0044) <= sig_slow(0043) or sig_fast(0150) or sig_slow(0029) or sig_slow(0022) or sig_slow(0013);
sig_slow(0045) <= sig_slow(0044) or sig_fast(0019) or sig_slow(0008) or sig_slow(0023) or sig_slow(0010);
sig_slow(0046) <= sig_slow(0045) or sig_fast(0015) or sig_slow(0037) or sig_slow(0026) or sig_slow(0000);
sig_slow(0047) <= sig_slow(0046) or sig_fast(0013) or sig_slow(0032) or sig_slow(0034) or sig_slow(0002);
sig_slow(0048) <= sig_slow(0047) or sig_fast(0050) or sig_slow(0047) or sig_slow(0032) or sig_slow(0023);
sig_slow(0049) <= sig_slow(0048) or sig_fast(0163) or sig_slow(0017) or sig_slow(0008) or sig_slow(0044);
sig_slow(0050) <= sig_slow(0049) or sig_fast(0126) or sig_slow(0034) or sig_slow(0010) or sig_slow(0036);
sig_slow(0051) <= sig_slow(0050) or sig_fast(0113) or sig_slow(0011) or sig_slow(0011) or sig_slow(0046);
sig_slow(0052) <= sig_slow(0051) or sig_fast(0052) or sig_slow(0042) or sig_slow(0024) or sig_slow(0010);
sig_slow(0053) <= sig_slow(0052) or sig_fast(0007) or sig_slow(0034) or sig_slow(0028) or sig_slow(0000);
sig_slow(0054) <= sig_slow(0053) or sig_fast(0044) or sig_slow(0016) or sig_slow(0024) or sig_slow(0004);
sig_slow(0055) <= sig_slow(0054) or sig_fast(0154) or sig_slow(0025) or sig_slow(0037) or sig_slow(0022);
sig_slow(0056) <= sig_slow(0055) or sig_fast(0140) or sig_slow(0013) or sig_slow(0031) or sig_slow(0013);
sig_slow(0057) <= sig_slow(0056) or sig_fast(0045) or sig_slow(0036) or sig_slow(0029) or sig_slow(0000);
sig_slow(0058) <= sig_slow(0057) or sig_fast(0000) or sig_slow(0052) or sig_slow(0000) or sig_slow(0011);
sig_slow(0059) <= sig_slow(0058) or sig_fast(0043) or sig_slow(0030) or sig_slow(0044) or sig_slow(0001);
sig_slow(0060) <= sig_slow(0059) or sig_fast(0122) or sig_slow(0008) or sig_slow(0007) or sig_slow(0024) or pushbutton;
sig_slow(0061) <= sig_slow(0060) or sig_fast(0144) or sig_slow(0038) or sig_slow(0046) or sig_slow(0029);
sig_slow(0062) <= sig_slow(0061) or sig_fast(0095) or sig_slow(0002) or sig_slow(0036) or sig_slow(0008);
sig_slow(0063) <= sig_slow(0062) or sig_fast(0089) or sig_slow(0034) or sig_slow(0052) or sig_slow(0018);
sig_slow(0064) <= sig_slow(0063) or sig_fast(0008) or sig_slow(0040) or sig_slow(0005) or sig_slow(0018);
sig_slow(0065) <= sig_slow(0064) or sig_fast(0103) or sig_slow(0017) or sig_slow(0019) or sig_slow(0002);
sig_slow(0066) <= sig_slow(0065) or sig_fast(0049) or sig_slow(0037) or sig_slow(0048) or sig_slow(0043);
sig_slow(0067) <= sig_slow(0066) or sig_fast(0005) or sig_slow(0063) or sig_slow(0002) or sig_slow(0029);
sig_slow(0068) <= sig_slow(0067) or sig_fast(0033) or sig_slow(0007) or sig_slow(0006) or sig_slow(0067);
sig_slow(0069) <= sig_slow(0068) or sig_fast(0005) or sig_slow(0067) or sig_slow(0003) or sig_slow(0067);
sig_slow(0070) <= sig_slow(0069) or sig_fast(0043) or sig_slow(0048) or sig_slow(0030) or sig_slow(0003);
sig_slow(0071) <= sig_slow(0070) or sig_fast(0155) or sig_slow(0042) or sig_slow(0058) or sig_slow(0037);
sig_slow(0072) <= sig_slow(0071) or sig_fast(0152) or sig_slow(0001) or sig_slow(0033) or sig_slow(0042);
sig_slow(0073) <= sig_slow(0072) or sig_fast(0116) or sig_slow(0031) or sig_slow(0066) or sig_slow(0015);
sig_slow(0074) <= sig_slow(0073) or sig_fast(0051) or sig_slow(0025) or sig_slow(0060) or sig_slow(0041);
sig_slow(0075) <= sig_slow(0074) or sig_fast(0073) or sig_slow(0023) or sig_slow(0017) or sig_slow(0027);
sig_slow(0076) <= sig_slow(0075) or sig_fast(0146) or sig_slow(0048) or sig_slow(0010) or sig_slow(0064);
sig_slow(0077) <= sig_slow(0076) or sig_fast(0066) or sig_slow(0051) or sig_slow(0024) or sig_slow(0010);
sig_slow(0078) <= sig_slow(0077) or sig_fast(0061) or sig_slow(0072) or sig_slow(0009) or sig_slow(0007);
sig_slow(0079) <= sig_slow(0078) or sig_fast(0129) or sig_slow(0023) or sig_slow(0004) or sig_slow(0073);
sig_slow(0080) <= sig_slow(0079) or sig_fast(0135) or sig_slow(0016) or sig_slow(0038) or sig_slow(0043) or pushbutton;
sig_slow(0081) <= sig_slow(0080) or sig_fast(0180) or sig_slow(0033) or sig_slow(0069) or sig_slow(0070);
sig_slow(0082) <= sig_slow(0081) or sig_fast(0000) or sig_slow(0080) or sig_slow(0073) or sig_slow(0021);
sig_slow(0083) <= sig_slow(0082) or sig_fast(0016) or sig_slow(0058) or sig_slow(0067) or sig_slow(0016);
sig_slow(0084) <= sig_slow(0083) or sig_fast(0172) or sig_slow(0006) or sig_slow(0027) or sig_slow(0065);
sig_slow(0085) <= sig_slow(0084) or sig_fast(0156) or sig_slow(0013) or sig_slow(0016) or sig_slow(0046);
sig_slow(0086) <= sig_slow(0085) or sig_fast(0040) or sig_slow(0040) or sig_slow(0060) or sig_slow(0053);
sig_slow(0087) <= sig_slow(0086) or sig_fast(0128) or sig_slow(0064) or sig_slow(0016) or sig_slow(0015);
sig_slow(0088) <= sig_slow(0087) or sig_fast(0046) or sig_slow(0049) or sig_slow(0034) or sig_slow(0065);
sig_slow(0089) <= sig_slow(0088) or sig_fast(0026) or sig_slow(0026) or sig_slow(0034) or sig_slow(0059);
sig_slow(0090) <= sig_slow(0089) or sig_fast(0079) or sig_slow(0066) or sig_slow(0079) or sig_slow(0001);
sig_slow(0091) <= sig_slow(0090) or sig_fast(0018) or sig_slow(0002) or sig_slow(0041) or sig_slow(0025);
sig_slow(0092) <= sig_slow(0091) or sig_fast(0094) or sig_slow(0073) or sig_slow(0028) or sig_slow(0043);
sig_slow(0093) <= sig_slow(0092) or sig_fast(0097) or sig_slow(0033) or sig_slow(0086) or sig_slow(0001);
sig_slow(0094) <= sig_slow(0093) or sig_fast(0186) or sig_slow(0065) or sig_slow(0015) or sig_slow(0062);
sig_slow(0095) <= sig_slow(0094) or sig_fast(0180) or sig_slow(0052) or sig_slow(0008) or sig_slow(0040);
sig_slow(0096) <= sig_slow(0095) or sig_fast(0098) or sig_slow(0014) or sig_slow(0038) or sig_slow(0067);
sig_slow(0097) <= sig_slow(0096) or sig_fast(0122) or sig_slow(0043) or sig_slow(0012) or sig_slow(0029);
sig_slow(0098) <= sig_slow(0097) or sig_fast(0121) or sig_slow(0005) or sig_slow(0070) or sig_slow(0082);
sig_slow(0099) <= sig_slow(0098) or sig_fast(0013) or sig_slow(0000) or sig_slow(0064) or sig_slow(0050);
sig_slow(0100) <= sig_slow(0099) or sig_fast(0177) or sig_slow(0081) or sig_slow(0051) or sig_slow(0088) or pushbutton;
sig_slow(0101) <= sig_slow(0100) or sig_fast(0183) or sig_slow(0024) or sig_slow(0055) or sig_slow(0055);
sig_slow(0102) <= sig_slow(0101) or sig_fast(0164) or sig_slow(0068) or sig_slow(0096) or sig_slow(0084);
sig_slow(0103) <= sig_slow(0102) or sig_fast(0044) or sig_slow(0072) or sig_slow(0092) or sig_slow(0011);
sig_slow(0104) <= sig_slow(0103) or sig_fast(0016) or sig_slow(0076) or sig_slow(0046) or sig_slow(0066);
sig_slow(0105) <= sig_slow(0104) or sig_fast(0118) or sig_slow(0010) or sig_slow(0003) or sig_slow(0001);
sig_slow(0106) <= sig_slow(0105) or sig_fast(0095) or sig_slow(0012) or sig_slow(0046) or sig_slow(0048);
sig_slow(0107) <= sig_slow(0106) or sig_fast(0150) or sig_slow(0105) or sig_slow(0036) or sig_slow(0006);
sig_slow(0108) <= sig_slow(0107) or sig_fast(0084) or sig_slow(0026) or sig_slow(0064) or sig_slow(0022);
sig_slow(0109) <= sig_slow(0108) or sig_fast(0089) or sig_slow(0072) or sig_slow(0049) or sig_slow(0019);
sig_slow(0110) <= sig_slow(0109) or sig_fast(0106) or sig_slow(0031) or sig_slow(0043) or sig_slow(0057);
sig_slow(0111) <= sig_slow(0110) or sig_fast(0062) or sig_slow(0074) or sig_slow(0110) or sig_slow(0082);
sig_slow(0112) <= sig_slow(0111) or sig_fast(0118) or sig_slow(0004) or sig_slow(0104) or sig_slow(0008);
sig_slow(0113) <= sig_slow(0112) or sig_fast(0096) or sig_slow(0093) or sig_slow(0043) or sig_slow(0037);
sig_slow(0114) <= sig_slow(0113) or sig_fast(0187) or sig_slow(0092) or sig_slow(0063) or sig_slow(0034);
sig_slow(0115) <= sig_slow(0114) or sig_fast(0195) or sig_slow(0114) or sig_slow(0001) or sig_slow(0074);
sig_slow(0116) <= sig_slow(0115) or sig_fast(0062) or sig_slow(0058) or sig_slow(0074) or sig_slow(0075);
sig_slow(0117) <= sig_slow(0116) or sig_fast(0163) or sig_slow(0021) or sig_slow(0008) or sig_slow(0075);
sig_slow(0118) <= sig_slow(0117) or sig_fast(0097) or sig_slow(0008) or sig_slow(0088) or sig_slow(0080);
sig_slow(0119) <= sig_slow(0118) or sig_fast(0174) or sig_slow(0011) or sig_slow(0092) or sig_slow(0083);
sig_slow(0120) <= sig_slow(0119) or sig_fast(0121) or sig_slow(0056) or sig_slow(0020) or sig_slow(0031) or pushbutton;
sig_slow(0121) <= sig_slow(0120) or sig_fast(0146) or sig_slow(0009) or sig_slow(0032) or sig_slow(0067);
sig_slow(0122) <= sig_slow(0121) or sig_fast(0162) or sig_slow(0043) or sig_slow(0047) or sig_slow(0032);
sig_slow(0123) <= sig_slow(0122) or sig_fast(0121) or sig_slow(0062) or sig_slow(0049) or sig_slow(0034);
sig_slow(0124) <= sig_slow(0123) or sig_fast(0091) or sig_slow(0105) or sig_slow(0050) or sig_slow(0105);
sig_slow(0125) <= sig_slow(0124) or sig_fast(0139) or sig_slow(0038) or sig_slow(0014) or sig_slow(0107);
sig_slow(0126) <= sig_slow(0125) or sig_fast(0036) or sig_slow(0049) or sig_slow(0100) or sig_slow(0009);
sig_slow(0127) <= sig_slow(0126) or sig_fast(0107) or sig_slow(0007) or sig_slow(0049) or sig_slow(0017);
sig_slow(0128) <= sig_slow(0127) or sig_fast(0173) or sig_slow(0089) or sig_slow(0005) or sig_slow(0072);
sig_slow(0129) <= sig_slow(0128) or sig_fast(0047) or sig_slow(0021) or sig_slow(0025) or sig_slow(0023);
sig_slow(0130) <= sig_slow(0129) or sig_fast(0136) or sig_slow(0061) or sig_slow(0087) or sig_slow(0089);
sig_slow(0131) <= sig_slow(0130) or sig_fast(0037) or sig_slow(0021) or sig_slow(0060) or sig_slow(0059);
sig_slow(0132) <= sig_slow(0131) or sig_fast(0115) or sig_slow(0012) or sig_slow(0096) or sig_slow(0130);
sig_slow(0133) <= sig_slow(0132) or sig_fast(0054) or sig_slow(0108) or sig_slow(0009) or sig_slow(0083);
sig_slow(0134) <= sig_slow(0133) or sig_fast(0175) or sig_slow(0101) or sig_slow(0117) or sig_slow(0103);
sig_slow(0135) <= sig_slow(0134) or sig_fast(0112) or sig_slow(0086) or sig_slow(0133) or sig_slow(0067);
sig_slow(0136) <= sig_slow(0135) or sig_fast(0057) or sig_slow(0033) or sig_slow(0116) or sig_slow(0000);
sig_slow(0137) <= sig_slow(0136) or sig_fast(0096) or sig_slow(0128) or sig_slow(0055) or sig_slow(0100);
sig_slow(0138) <= sig_slow(0137) or sig_fast(0126) or sig_slow(0078) or sig_slow(0088) or sig_slow(0015);
sig_slow(0139) <= sig_slow(0138) or sig_fast(0146) or sig_slow(0039) or sig_slow(0034) or sig_slow(0047);
sig_slow(0140) <= sig_slow(0139) or sig_fast(0199) or sig_slow(0137) or sig_slow(0064) or sig_slow(0058) or pushbutton;
sig_slow(0141) <= sig_slow(0140) or sig_fast(0013) or sig_slow(0059) or sig_slow(0032) or sig_slow(0038);
sig_slow(0142) <= sig_slow(0141) or sig_fast(0123) or sig_slow(0094) or sig_slow(0112) or sig_slow(0077);
sig_slow(0143) <= sig_slow(0142) or sig_fast(0051) or sig_slow(0101) or sig_slow(0034) or sig_slow(0100);
sig_slow(0144) <= sig_slow(0143) or sig_fast(0152) or sig_slow(0034) or sig_slow(0006) or sig_slow(0061);
sig_slow(0145) <= sig_slow(0144) or sig_fast(0100) or sig_slow(0030) or sig_slow(0118) or sig_slow(0117);
sig_slow(0146) <= sig_slow(0145) or sig_fast(0154) or sig_slow(0122) or sig_slow(0143) or sig_slow(0059);
sig_slow(0147) <= sig_slow(0146) or sig_fast(0109) or sig_slow(0137) or sig_slow(0002) or sig_slow(0053);
sig_slow(0148) <= sig_slow(0147) or sig_fast(0169) or sig_slow(0121) or sig_slow(0114) or sig_slow(0059);
sig_slow(0149) <= sig_slow(0148) or sig_fast(0142) or sig_slow(0135) or sig_slow(0144) or sig_slow(0053);
sig_slow(0150) <= sig_slow(0149) or sig_fast(0141) or sig_slow(0052) or sig_slow(0136) or sig_slow(0008);
sig_slow(0151) <= sig_slow(0150) or sig_fast(0102) or sig_slow(0048) or sig_slow(0141) or sig_slow(0044);
sig_slow(0152) <= sig_slow(0151) or sig_fast(0098) or sig_slow(0139) or sig_slow(0090) or sig_slow(0010);
sig_slow(0153) <= sig_slow(0152) or sig_fast(0099) or sig_slow(0074) or sig_slow(0091) or sig_slow(0034);
sig_slow(0154) <= sig_slow(0153) or sig_fast(0171) or sig_slow(0006) or sig_slow(0072) or sig_slow(0150);
sig_slow(0155) <= sig_slow(0154) or sig_fast(0111) or sig_slow(0020) or sig_slow(0022) or sig_slow(0040);
sig_slow(0156) <= sig_slow(0155) or sig_fast(0033) or sig_slow(0131) or sig_slow(0127) or sig_slow(0061);
sig_slow(0157) <= sig_slow(0156) or sig_fast(0008) or sig_slow(0111) or sig_slow(0047) or sig_slow(0018);
sig_slow(0158) <= sig_slow(0157) or sig_fast(0131) or sig_slow(0056) or sig_slow(0155) or sig_slow(0060);
sig_slow(0159) <= sig_slow(0158) or sig_fast(0050) or sig_slow(0035) or sig_slow(0031) or sig_slow(0030);
sig_slow(0160) <= sig_slow(0159) or sig_fast(0100) or sig_slow(0131) or sig_slow(0032) or sig_slow(0098) or pushbutton;
sig_slow(0161) <= sig_slow(0160) or sig_fast(0027) or sig_slow(0146) or sig_slow(0067) or sig_slow(0092);
sig_slow(0162) <= sig_slow(0161) or sig_fast(0087) or sig_slow(0149) or sig_slow(0017) or sig_slow(0063);
sig_slow(0163) <= sig_slow(0162) or sig_fast(0103) or sig_slow(0029) or sig_slow(0040) or sig_slow(0131);
sig_slow(0164) <= sig_slow(0163) or sig_fast(0045) or sig_slow(0094) or sig_slow(0096) or sig_slow(0051);
sig_slow(0165) <= sig_slow(0164) or sig_fast(0129) or sig_slow(0116) or sig_slow(0097) or sig_slow(0156);
sig_slow(0166) <= sig_slow(0165) or sig_fast(0008) or sig_slow(0100) or sig_slow(0162) or sig_slow(0031);
sig_slow(0167) <= sig_slow(0166) or sig_fast(0089) or sig_slow(0028) or sig_slow(0059) or sig_slow(0106);
sig_slow(0168) <= sig_slow(0167) or sig_fast(0171) or sig_slow(0134) or sig_slow(0098) or sig_slow(0005);
sig_slow(0169) <= sig_slow(0168) or sig_fast(0074) or sig_slow(0054) or sig_slow(0158) or sig_slow(0128);
sig_slow(0170) <= sig_slow(0169) or sig_fast(0177) or sig_slow(0092) or sig_slow(0023) or sig_slow(0048);
sig_slow(0171) <= sig_slow(0170) or sig_fast(0178) or sig_slow(0092) or sig_slow(0108) or sig_slow(0063);
sig_slow(0172) <= sig_slow(0171) or sig_fast(0019) or sig_slow(0118) or sig_slow(0062) or sig_slow(0163);
sig_slow(0173) <= sig_slow(0172) or sig_fast(0067) or sig_slow(0134) or sig_slow(0041) or sig_slow(0158);
sig_slow(0174) <= sig_slow(0173) or sig_fast(0162) or sig_slow(0101) or sig_slow(0044) or sig_slow(0133);
sig_slow(0175) <= sig_slow(0174) or sig_fast(0079) or sig_slow(0137) or sig_slow(0027) or sig_slow(0106);
sig_slow(0176) <= sig_slow(0175) or sig_fast(0050) or sig_slow(0138) or sig_slow(0158) or sig_slow(0028);
sig_slow(0177) <= sig_slow(0176) or sig_fast(0148) or sig_slow(0141) or sig_slow(0009) or sig_slow(0102);
sig_slow(0178) <= sig_slow(0177) or sig_fast(0060) or sig_slow(0079) or sig_slow(0060) or sig_slow(0025);
sig_slow(0179) <= sig_slow(0178) or sig_fast(0069) or sig_slow(0108) or sig_slow(0080) or sig_slow(0148);
sig_slow(0180) <= sig_slow(0179) or sig_fast(0140) or sig_slow(0101) or sig_slow(0036) or sig_slow(0059) or pushbutton;
sig_slow(0181) <= sig_slow(0180) or sig_fast(0026) or sig_slow(0161) or sig_slow(0170) or sig_slow(0137);
sig_slow(0182) <= sig_slow(0181) or sig_fast(0018) or sig_slow(0035) or sig_slow(0049) or sig_slow(0097);
sig_slow(0183) <= sig_slow(0182) or sig_fast(0185) or sig_slow(0006) or sig_slow(0026) or sig_slow(0000);
sig_slow(0184) <= sig_slow(0183) or sig_fast(0174) or sig_slow(0053) or sig_slow(0127) or sig_slow(0098);
sig_slow(0185) <= sig_slow(0184) or sig_fast(0182) or sig_slow(0115) or sig_slow(0090) or sig_slow(0141);
sig_slow(0186) <= sig_slow(0185) or sig_fast(0052) or sig_slow(0034) or sig_slow(0011) or sig_slow(0120);
sig_slow(0187) <= sig_slow(0186) or sig_fast(0007) or sig_slow(0142) or sig_slow(0063) or sig_slow(0092);
sig_slow(0188) <= sig_slow(0187) or sig_fast(0124) or sig_slow(0065) or sig_slow(0145) or sig_slow(0064);
sig_slow(0189) <= sig_slow(0188) or sig_fast(0090) or sig_slow(0100) or sig_slow(0141) or sig_slow(0118);
sig_slow(0190) <= sig_slow(0189) or sig_fast(0011) or sig_slow(0109) or sig_slow(0109) or sig_slow(0163);
sig_slow(0191) <= sig_slow(0190) or sig_fast(0147) or sig_slow(0045) or sig_slow(0115) or sig_slow(0125);
sig_slow(0192) <= sig_slow(0191) or sig_fast(0147) or sig_slow(0004) or sig_slow(0181) or sig_slow(0105);
sig_slow(0193) <= sig_slow(0192) or sig_fast(0132) or sig_slow(0124) or sig_slow(0046) or sig_slow(0170);
sig_slow(0194) <= sig_slow(0193) or sig_fast(0194) or sig_slow(0148) or sig_slow(0090) or sig_slow(0039);
sig_slow(0195) <= sig_slow(0194) or sig_fast(0110) or sig_slow(0162) or sig_slow(0189) or sig_slow(0179);
sig_slow(0196) <= sig_slow(0195) or sig_fast(0195) or sig_slow(0046) or sig_slow(0114) or sig_slow(0022);
sig_slow(0197) <= sig_slow(0196) or sig_fast(0156) or sig_slow(0174) or sig_slow(0189) or sig_slow(0073);
sig_slow(0198) <= sig_slow(0197) or sig_fast(0087) or sig_slow(0177) or sig_slow(0170) or sig_slow(0064);
sig_slow(0199) <= sig_slow(0198) or sig_fast(0090) or sig_slow(0022) or sig_slow(0171) or sig_slow(0194);
reset_global <= sig_slow(0) or sig_slow(0000) or sig_slow(0020) or sig_slow(0040) or sig_slow(0060) or sig_slow(0080) or sig_slow(0100) or sig_slow(0120) or sig_slow(0140) or sig_slow(0160) or sig_slow(0180) or sig_slow(0200);
                
        end if;
end process;

end rst_mgr_arch;


